module robot ( 
	a,
	b,
	c,
	d,
	e,
	f1,
	f2
	) ;

input  a;
input  b;
input  c;
input  d;
input  e;
inout  f1;
inout  f2;
