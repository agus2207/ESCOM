module det ( 
	en,
	clk,
	clr,
	s
	) ;

input  en;
input  clk;
input  clr;
inout  s;
