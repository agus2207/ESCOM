module suma ( 
	a,
	b,
	control,
	clk,
	clr,
	c,
	s
	) ;

input  a;
input  b;
input  control;
input  clk;
input  clr;
inout  c;
inout [3:0] s;
