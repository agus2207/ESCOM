module det ( 
	en,
	clk,
	s
	) ;

input  en;
input  clk;
inout  s;
